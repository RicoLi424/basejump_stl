/**
 *    bsg_cache_dma_to_wormhole.v
 *
 *    This module interfaces bsg_cache_nb_dma to a wormhole link.
 *    dma_pkts come in two flavors:
 *      - Write packets send a wormhole header flit, then an address flit, a mask flit, then N data flits (the
 *          evicted data)
 *      - Read packets send a wormhole header flit, then an address flit, an mshr id flit, then receive
 *          N data flits (the fill data) and mshr id flit asynchronously.
 */

`include "bsg_defines.v"
`include "bsg_noc_links.vh"
`include "bsg_cache_nb.vh"

module bsg_cache_nb_dma_to_wormhole
 import bsg_noc_pkg::*;
 import bsg_cache_nb_pkg::*;
 #(parameter `BSG_INV_PARAM(dma_addr_width_p) // cache addr width (byte addr)
   , parameter `BSG_INV_PARAM(block_size_in_bursts_p) // num of data beats in dma transfer
   , parameter `BSG_INV_PARAM(dma_mask_width_p) // mask width in the bsg_cache_dma_pkt_s. This should equal to the block_size_in_words_p set for bsg_cache_nb.

   , parameter `BSG_INV_PARAM(mshr_els_p)

   // flit width should match the cache dma width.
   , parameter `BSG_INV_PARAM(wh_flit_width_p)
   , parameter `BSG_INV_PARAM(wh_cid_width_p)
   , parameter `BSG_INV_PARAM(wh_len_width_p)
   , parameter `BSG_INV_PARAM(wh_cord_width_p)

   , parameter dma_pkt_width_lp=`bsg_cache_nb_dma_pkt_width(dma_addr_width_p, dma_mask_width_p, mshr_els_p)
   , parameter wh_link_sif_width_lp=`bsg_ready_and_link_sif_width(wh_flit_width_p)
   , parameter dma_data_width_lp=wh_flit_width_p

   , parameter lg_mshr_els_lp = `BSG_SAFE_CLOG2(mshr_els_p)

   // Whether to buffer the returning data flits. May be necessary for timing purposes
   , parameter buffer_return_p = 1
   )
  (
   input clk_i
   , input reset_i

   , input [dma_pkt_width_lp-1:0] dma_pkt_i
   , input dma_pkt_v_i
   , output dma_pkt_yumi_o

   , output logic [dma_data_width_lp-1:0] dma_data_o
   , output logic [lg_mshr_els_lp-1:0] dma_mshr_id_o
   , output logic dma_data_v_o
   , input dma_data_ready_and_i

   , input [dma_data_width_lp-1:0] dma_data_i
   , input dma_data_v_i
   , output logic dma_data_yumi_o

   , input [wh_link_sif_width_lp-1:0] wh_link_sif_i
   , output logic [wh_link_sif_width_lp-1:0] wh_link_sif_o

   , input [wh_cord_width_p-1:0] my_wh_cord_i
   , input [wh_cord_width_p-1:0] dest_wh_cord_i
   , input [wh_cid_width_p-1:0] my_wh_cid_i
   , input [wh_cid_width_p-1:0] dest_wh_cid_i
   );

  `declare_bsg_cache_nb_dma_pkt_s(dma_addr_width_p, dma_mask_width_p, mshr_els_p);
  `declare_bsg_ready_and_link_sif_s(wh_flit_width_p, wh_link_sif_s);
  wh_link_sif_s wh_link_sif_in;
  wh_link_sif_s wh_link_sif_out;
  assign wh_link_sif_in = wh_link_sif_i;
  assign wh_link_sif_o = wh_link_sif_out;

  // dma pkt fifo
  logic dma_pkt_ready_lo;
  logic dma_pkt_v_lo;
  logic dma_pkt_yumi_li;
  bsg_cache_nb_dma_pkt_s dma_pkt_lo;


  bsg_fifo_1r1w_small #(
    .width_p(dma_pkt_width_lp)
    ,.els_p(mshr_els_p*2)
  ) dma_pkt_fifo (
    .clk_i(clk_i)
    ,.reset_i(reset_i)
    ,.data_i(dma_pkt_i)
    ,.v_i(dma_pkt_v_i)
    ,.ready_o(dma_pkt_ready_lo)
    ,.v_o(dma_pkt_v_lo)
    ,.data_o(dma_pkt_lo)
    ,.yumi_i(dma_pkt_yumi_li)
  );

  assign dma_pkt_yumi_o = dma_pkt_ready_lo & dma_pkt_v_i;


  logic evict_data_fifo_ready_lo;
  logic evict_data_fifo_v_lo, evict_data_fifo_yumi_li;
  logic [dma_data_width_lp-1:0] evict_data_fifo_data_lo;

  bsg_fifo_1r1w_small #(
    .width_p(wh_flit_width_p)
    ,.els_p(mshr_els_p*block_size_in_bursts_p)
  ) evict_data_fifo (
    .clk_i      (clk_i)
    ,.reset_i   (reset_i)

    ,.v_i       (dma_data_v_i)
    ,.data_i    (dma_data_i)
    ,.ready_o   (evict_data_fifo_ready_lo)

    ,.v_o       (evict_data_fifo_v_lo)
    ,.data_o    (evict_data_fifo_data_lo)
    ,.yumi_i    (evict_data_fifo_yumi_li)
  );

  assign dma_data_yumi_o = evict_data_fifo_ready_lo & dma_data_v_i;


  // FIFO for wormhole flits coming back to vcache.
  logic return_data_fifo_v_lo;
  logic [wh_flit_width_p-1:0] return_data_fifo_data_lo;
  logic return_data_fifo_ready_li, return_data_fifo_yumi_li;

  if (buffer_return_p) begin : br
    bsg_fifo_1r1w_small #(
      .width_p(wh_flit_width_p)
      ,.els_p(mshr_els_p*(1+block_size_in_bursts_p))
    ) return_data_fifo (
      .clk_i      (clk_i)
      ,.reset_i   (reset_i)

      ,.v_i       (wh_link_sif_in.v)
      ,.data_i    (wh_link_sif_in.data)
      ,.ready_o   (wh_link_sif_out.ready_and_rev)

      ,.v_o       (return_data_fifo_v_lo)
      ,.data_o    (return_data_fifo_data_lo)
      ,.yumi_i    (return_data_fifo_yumi_li)
    );
    assign return_data_fifo_yumi_li = return_data_fifo_ready_li & return_data_fifo_v_lo;


  end else begin : nbr
    assign return_data_fifo_v_lo = wh_link_sif_in.v;
    assign return_data_fifo_data_lo = wh_link_sif_in.data;
    assign wh_link_sif_out.ready_and_rev = return_data_fifo_ready_li;
    assign return_data_fifo_yumi_li = wh_link_sif_out.ready_and_rev & wh_link_sif_in.v;
  end


  // counter
  localparam count_width_lp = `BSG_SAFE_CLOG2(block_size_in_bursts_p);
  logic send_clear_li;
  logic send_up_li;
  logic [count_width_lp-1:0] send_count_lo;

  bsg_counter_clear_up #(
    .max_val_p(block_size_in_bursts_p-1)
    ,.init_val_p(0)
  ) send_count (
    .clk_i(clk_i)
    ,.reset_i(reset_i)
    ,.clear_i(send_clear_li)
    ,.up_i(send_up_li)
    ,.count_o(send_count_lo)
  );

  // send FSM
  enum logic [2:0] {
    SEND_RESET
    , SEND_READY
    , SEND_ADDR
    , SEND_MASK
    , SEND_DATA
  } send_state_n, send_state_r;


  // Check if mask bits are all 1.
  wire mask_all_one = &dma_pkt_lo.mask;

  // Make a header flit.
  `declare_bsg_cache_nb_wh_header_flit_s(wh_flit_width_p,wh_cord_width_p,wh_len_width_p,wh_cid_width_p,mshr_els_p);

  bsg_cache_nb_wh_header_flit_s send_header_flit;
  assign send_header_flit.unused = '0;
  assign send_header_flit.opcode = dma_pkt_lo.write_not_read
    ? (mask_all_one 
      ? e_cache_wh_write_non_masked 
      : e_cache_wh_write_masked)
    : e_cache_wh_read;
  assign send_header_flit.mshr_id = dma_pkt_lo.mshr_id;
  assign send_header_flit.src_cid = my_wh_cid_i;
  assign send_header_flit.src_cord = my_wh_cord_i;
  assign send_header_flit.len = dma_pkt_lo.write_not_read
    ? (mask_all_one 
      ? wh_len_width_p'(1+block_size_in_bursts_p) // header + addr + data
      : wh_len_width_p'(2+block_size_in_bursts_p)) // header + addr + mask + data
    : wh_len_width_p'(1);  // header + addr
  assign send_header_flit.cord = dest_wh_cord_i;
  assign send_header_flit.cid = dest_wh_cid_i;


  always_comb begin

    send_state_n = send_state_r;
    dma_pkt_yumi_li = 1'b0;
    send_clear_li = 1'b0;
    send_up_li = 1'b0;
    wh_link_sif_out.v = 1'b0;
    wh_link_sif_out.data = evict_data_fifo_data_lo;
    evict_data_fifo_yumi_li = 1'b0;

    case (send_state_r)
      SEND_RESET: begin
        send_state_n = SEND_READY;
      end

      SEND_READY: begin
        // send header
        wh_link_sif_out.data = send_header_flit;
        if (dma_pkt_v_lo) begin
          wh_link_sif_out.v = 1'b1;
          send_state_n = (wh_link_sif_in.ready_and_rev)
            ? SEND_ADDR
            : SEND_READY;
        end
      end

      SEND_ADDR: begin
        wh_link_sif_out.data = wh_flit_width_p'(dma_pkt_lo.addr);
        if (dma_pkt_v_lo) begin
          wh_link_sif_out.v = 1'b1;
 
          // If it's read, dequeue dma_pkt.
          // If it's masked write, don't dequeue yet, because it still needs to send the mask flit.
          // If it's non-masked write, dequeue it .
          dma_pkt_yumi_li = dma_pkt_lo.write_not_read
            ? (mask_all_one
              ? wh_link_sif_in.ready_and_rev  // non-masked write
              : 1'b0)  // masked write
            : wh_link_sif_in.ready_and_rev;

          send_state_n = wh_link_sif_in.ready_and_rev
            ? (dma_pkt_lo.write_not_read 
              ? (mask_all_one ? SEND_DATA : SEND_MASK)
              : SEND_READY)
            : SEND_ADDR;
        end
      end
    
      SEND_MASK: begin
        wh_link_sif_out.data = wh_flit_width_p'(dma_pkt_lo.mask);
        if (dma_pkt_v_lo) begin
          wh_link_sif_out.v = 1'b1;
          dma_pkt_yumi_li = wh_link_sif_in.ready_and_rev;
          send_state_n = wh_link_sif_in.ready_and_rev
            ? SEND_DATA
            : SEND_MASK;
        end
      end

      SEND_DATA: begin
        wh_link_sif_out.data = evict_data_fifo_data_lo;
        if (evict_data_fifo_v_lo) begin
          wh_link_sif_out.v = 1'b1;
          evict_data_fifo_yumi_li = wh_link_sif_in.ready_and_rev & wh_link_sif_out.v;
          send_up_li = evict_data_fifo_yumi_li & (send_count_lo != block_size_in_bursts_p-1);
          send_clear_li = evict_data_fifo_yumi_li & (send_count_lo == block_size_in_bursts_p-1);
          send_state_n = send_clear_li
            ? SEND_READY
            : SEND_DATA;
        end
      end

      // should never happen
      default: begin
        send_state_n = SEND_READY;
      end
    endcase
  end

  bsg_cache_nb_wh_header_flit_s return_header_flit;
  assign return_header_flit = return_data_fifo_data_lo;

  // receiver FSM
  logic recv_clear_li;
  logic recv_up_li;
  logic [count_width_lp-1:0] recv_count_lo;

  bsg_counter_clear_up #(
    .max_val_p(block_size_in_bursts_p-1)
    ,.init_val_p(0)
  ) recv_count (
    .clk_i(clk_i)
    ,.reset_i(reset_i)
    ,.clear_i(recv_clear_li)
    ,.up_i(recv_up_li)
    ,.count_o(recv_count_lo)
  );

  typedef enum logic [1:0] {
    RECV_RESET
    , RECV_READY
    , RECV_DATA
  } recv_state_e;

  recv_state_e recv_state_r, recv_state_n;

  logic [lg_mshr_els_lp-1:0] refill_mshr_id_r, refill_mshr_id_n;

  always_comb begin
    recv_state_n = recv_state_r;
    recv_clear_li = 1'b0;
    recv_up_li = 1'b0;
    return_data_fifo_ready_li = 1'b0;
    dma_data_v_o = 1'b0;
    dma_data_o = return_data_fifo_data_lo;
    dma_mshr_id_o = refill_mshr_id_r;
    refill_mshr_id_n = refill_mshr_id_r;

    case (recv_state_r)
      RECV_RESET: begin
        recv_state_n = RECV_READY;
      end

      RECV_READY: begin
        return_data_fifo_ready_li = 1'b1;
        refill_mshr_id_n = return_data_fifo_yumi_li ? return_header_flit.mshr_id : refill_mshr_id_r;
        recv_state_n = return_data_fifo_yumi_li
          ? RECV_DATA
          : RECV_READY;
      end

      RECV_DATA: begin
        return_data_fifo_ready_li = dma_data_ready_and_i;
        dma_data_v_o = return_data_fifo_v_lo;
        recv_up_li = return_data_fifo_yumi_li & (recv_count_lo != block_size_in_bursts_p-1);
        recv_clear_li = return_data_fifo_yumi_li & (recv_count_lo == block_size_in_bursts_p-1);
        recv_state_n = recv_clear_li
          ? RECV_READY
          : RECV_DATA;
      end

      default: begin
        recv_state_n = RECV_READY;
      end
    endcase
  end




  // sequential logic
  // synopsys sync_set_reset "reset_i"
  always_ff @ (posedge clk_i) begin
    if (reset_i) begin
      send_state_r <= SEND_RESET;
      recv_state_r <= RECV_RESET;
      refill_mshr_id_r <= '0;
    end
    else begin
      send_state_r <= send_state_n;
      recv_state_r <= recv_state_n;
      refill_mshr_id_r <= refill_mshr_id_n;
    end
  end

  //synopsys translate_off
  if (wh_flit_width_p != dma_data_width_lp)
    $error("WH flit width must be equal to DMA data width");
  if (wh_flit_width_p < dma_addr_width_p)
    $error("WH flit width must be larger than address width");
  if (wh_len_width_p < `BSG_WIDTH(block_size_in_bursts_p+1))
    $error("WH len width %d must be large enough to hold the dma transfer size %d", wh_len_width_p, `BSG_WIDTH(block_size_in_bursts_p+1));
  //synopsys translate_on

endmodule

`BSG_ABSTRACT_MODULE(bsg_cache_nb_dma_to_wormhole)
